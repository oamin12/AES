module ShiftRows_tb();

reg [127:0] inputValue;
wire [127:0] outputValue;


initial begin 
 $monitor ("%h   %h", 
  	  inputValue, outputValue);
	  
inputValue = 127'h 63cab7040953d051cd60e0e7ba70e18c;



end
ShiftRows v(inputValue, outputValue);


endmodule 