module sbox(input wire [31 : 0]  inputSbox,output wire [31 : 0] outputSbox);


  wire [7 : 0] lookUpTable [0 : 255];



  assign outputSbox[31 : 24] = lookUpTable[inputSbox[31 : 24]];
  assign outputSbox[23 : 16] = lookUpTable[inputSbox[23 : 16]];
  assign outputSbox[15 : 08] = lookUpTable[inputSbox[15 : 08]];
  assign outputSbox[07 : 00] = lookUpTable[inputSbox[07 : 00]];


  assign lookUpTable[8'h00] = 8'h63;
  assign lookUpTable[8'h01] = 8'h7c;
  assign lookUpTable[8'h02] = 8'h77;
  assign lookUpTable[8'h03] = 8'h7b;
  assign lookUpTable[8'h04] = 8'hf2;
  assign lookUpTable[8'h05] = 8'h6b;
  assign lookUpTable[8'h06] = 8'h6f;
  assign lookUpTable[8'h07] = 8'hc5;
  assign lookUpTable[8'h08] = 8'h30;
  assign lookUpTable[8'h09] = 8'h01;
  assign lookUpTable[8'h0a] = 8'h67;
  assign lookUpTable[8'h0b] = 8'h2b;
  assign lookUpTable[8'h0c] = 8'hfe;
  assign lookUpTable[8'h0d] = 8'hd7;
  assign lookUpTable[8'h0e] = 8'hab;
  assign lookUpTable[8'h0f] = 8'h76;
  assign lookUpTable[8'h10] = 8'hca;
  assign lookUpTable[8'h11] = 8'h82;
  assign lookUpTable[8'h12] = 8'hc9;
  assign lookUpTable[8'h13] = 8'h7d;
  assign lookUpTable[8'h14] = 8'hfa;
  assign lookUpTable[8'h15] = 8'h59;
  assign lookUpTable[8'h16] = 8'h47;
  assign lookUpTable[8'h17] = 8'hf0;
  assign lookUpTable[8'h18] = 8'had;
  assign lookUpTable[8'h19] = 8'hd4;
  assign lookUpTable[8'h1a] = 8'ha2;
  assign lookUpTable[8'h1b] = 8'haf;
  assign lookUpTable[8'h1c] = 8'h9c;
  assign lookUpTable[8'h1d] = 8'ha4;
  assign lookUpTable[8'h1e] = 8'h72;
  assign lookUpTable[8'h1f] = 8'hc0;
  assign lookUpTable[8'h20] = 8'hb7;
  assign lookUpTable[8'h21] = 8'hfd;
  assign lookUpTable[8'h22] = 8'h93;
  assign lookUpTable[8'h23] = 8'h26;
  assign lookUpTable[8'h24] = 8'h36;
  assign lookUpTable[8'h25] = 8'h3f;
  assign lookUpTable[8'h26] = 8'hf7;
  assign lookUpTable[8'h27] = 8'hcc;
  assign lookUpTable[8'h28] = 8'h34;
  assign lookUpTable[8'h29] = 8'ha5;
  assign lookUpTable[8'h2a] = 8'he5;
  assign lookUpTable[8'h2b] = 8'hf1;
  assign lookUpTable[8'h2c] = 8'h71;
  assign lookUpTable[8'h2d] = 8'hd8;
  assign lookUpTable[8'h2e] = 8'h31;
  assign lookUpTable[8'h2f] = 8'h15;
  assign lookUpTable[8'h30] = 8'h04;
  assign lookUpTable[8'h31] = 8'hc7;
  assign lookUpTable[8'h32] = 8'h23;
  assign lookUpTable[8'h33] = 8'hc3;
  assign lookUpTable[8'h34] = 8'h18;
  assign lookUpTable[8'h35] = 8'h96;
  assign lookUpTable[8'h36] = 8'h05;
  assign lookUpTable[8'h37] = 8'h9a;
  assign lookUpTable[8'h38] = 8'h07;
  assign lookUpTable[8'h39] = 8'h12;
  assign lookUpTable[8'h3a] = 8'h80;
  assign lookUpTable[8'h3b] = 8'he2;
  assign lookUpTable[8'h3c] = 8'heb;
  assign lookUpTable[8'h3d] = 8'h27;
  assign lookUpTable[8'h3e] = 8'hb2;
  assign lookUpTable[8'h3f] = 8'h75;
  assign lookUpTable[8'h40] = 8'h09;
  assign lookUpTable[8'h41] = 8'h83;
  assign lookUpTable[8'h42] = 8'h2c;
  assign lookUpTable[8'h43] = 8'h1a;
  assign lookUpTable[8'h44] = 8'h1b;
  assign lookUpTable[8'h45] = 8'h6e;
  assign lookUpTable[8'h46] = 8'h5a;
  assign lookUpTable[8'h47] = 8'ha0;
  assign lookUpTable[8'h48] = 8'h52;
  assign lookUpTable[8'h49] = 8'h3b;
  assign lookUpTable[8'h4a] = 8'hd6;
  assign lookUpTable[8'h4b] = 8'hb3;
  assign lookUpTable[8'h4c] = 8'h29;
  assign lookUpTable[8'h4d] = 8'he3;
  assign lookUpTable[8'h4e] = 8'h2f;
  assign lookUpTable[8'h4f] = 8'h84;
  assign lookUpTable[8'h50] = 8'h53;
  assign lookUpTable[8'h51] = 8'hd1;
  assign lookUpTable[8'h52] = 8'h00;
  assign lookUpTable[8'h53] = 8'hed;
  assign lookUpTable[8'h54] = 8'h20;
  assign lookUpTable[8'h55] = 8'hfc;
  assign lookUpTable[8'h56] = 8'hb1;
  assign lookUpTable[8'h57] = 8'h5b;
  assign lookUpTable[8'h58] = 8'h6a;
  assign lookUpTable[8'h59] = 8'hcb;
  assign lookUpTable[8'h5a] = 8'hbe;
  assign lookUpTable[8'h5b] = 8'h39;
  assign lookUpTable[8'h5c] = 8'h4a;
  assign lookUpTable[8'h5d] = 8'h4c;
  assign lookUpTable[8'h5e] = 8'h58;
  assign lookUpTable[8'h5f] = 8'hcf;
  assign lookUpTable[8'h60] = 8'hd0;
  assign lookUpTable[8'h61] = 8'hef;
  assign lookUpTable[8'h62] = 8'haa;
  assign lookUpTable[8'h63] = 8'hfb;
  assign lookUpTable[8'h64] = 8'h43;
  assign lookUpTable[8'h65] = 8'h4d;
  assign lookUpTable[8'h66] = 8'h33;
  assign lookUpTable[8'h67] = 8'h85;
  assign lookUpTable[8'h68] = 8'h45;
  assign lookUpTable[8'h69] = 8'hf9;
  assign lookUpTable[8'h6a] = 8'h02;
  assign lookUpTable[8'h6b] = 8'h7f;
  assign lookUpTable[8'h6c] = 8'h50;
  assign lookUpTable[8'h6d] = 8'h3c;
  assign lookUpTable[8'h6e] = 8'h9f;
  assign lookUpTable[8'h6f] = 8'ha8;
  assign lookUpTable[8'h70] = 8'h51;
  assign lookUpTable[8'h71] = 8'ha3;
  assign lookUpTable[8'h72] = 8'h40;
  assign lookUpTable[8'h73] = 8'h8f;
  assign lookUpTable[8'h74] = 8'h92;
  assign lookUpTable[8'h75] = 8'h9d;
  assign lookUpTable[8'h76] = 8'h38;
  assign lookUpTable[8'h77] = 8'hf5;
  assign lookUpTable[8'h78] = 8'hbc;
  assign lookUpTable[8'h79] = 8'hb6;
  assign lookUpTable[8'h7a] = 8'hda;
  assign lookUpTable[8'h7b] = 8'h21;
  assign lookUpTable[8'h7c] = 8'h10;
  assign lookUpTable[8'h7d] = 8'hff;
  assign lookUpTable[8'h7e] = 8'hf3;
  assign lookUpTable[8'h7f] = 8'hd2;
  assign lookUpTable[8'h80] = 8'hcd;
  assign lookUpTable[8'h81] = 8'h0c;
  assign lookUpTable[8'h82] = 8'h13;
  assign lookUpTable[8'h83] = 8'hec;
  assign lookUpTable[8'h84] = 8'h5f;
  assign lookUpTable[8'h85] = 8'h97;
  assign lookUpTable[8'h86] = 8'h44;
  assign lookUpTable[8'h87] = 8'h17;
  assign lookUpTable[8'h88] = 8'hc4;
  assign lookUpTable[8'h89] = 8'ha7;
  assign lookUpTable[8'h8a] = 8'h7e;
  assign lookUpTable[8'h8b] = 8'h3d;
  assign lookUpTable[8'h8c] = 8'h64;
  assign lookUpTable[8'h8d] = 8'h5d;
  assign lookUpTable[8'h8e] = 8'h19;
  assign lookUpTable[8'h8f] = 8'h73;
  assign lookUpTable[8'h90] = 8'h60;
  assign lookUpTable[8'h91] = 8'h81;
  assign lookUpTable[8'h92] = 8'h4f;
  assign lookUpTable[8'h93] = 8'hdc;
  assign lookUpTable[8'h94] = 8'h22;
  assign lookUpTable[8'h95] = 8'h2a;
  assign lookUpTable[8'h96] = 8'h90;
  assign lookUpTable[8'h97] = 8'h88;
  assign lookUpTable[8'h98] = 8'h46;
  assign lookUpTable[8'h99] = 8'hee;
  assign lookUpTable[8'h9a] = 8'hb8;
  assign lookUpTable[8'h9b] = 8'h14;
  assign lookUpTable[8'h9c] = 8'hde;
  assign lookUpTable[8'h9d] = 8'h5e;
  assign lookUpTable[8'h9e] = 8'h0b;
  assign lookUpTable[8'h9f] = 8'hdb;
  assign lookUpTable[8'ha0] = 8'he0;
  assign lookUpTable[8'ha1] = 8'h32;
  assign lookUpTable[8'ha2] = 8'h3a;
  assign lookUpTable[8'ha3] = 8'h0a;
  assign lookUpTable[8'ha4] = 8'h49;
  assign lookUpTable[8'ha5] = 8'h06;
  assign lookUpTable[8'ha6] = 8'h24;
  assign lookUpTable[8'ha7] = 8'h5c;
  assign lookUpTable[8'ha8] = 8'hc2;
  assign lookUpTable[8'ha9] = 8'hd3;
  assign lookUpTable[8'haa] = 8'hac;
  assign lookUpTable[8'hab] = 8'h62;
  assign lookUpTable[8'hac] = 8'h91;
  assign lookUpTable[8'had] = 8'h95;
  assign lookUpTable[8'hae] = 8'he4;
  assign lookUpTable[8'haf] = 8'h79;
  assign lookUpTable[8'hb0] = 8'he7;
  assign lookUpTable[8'hb1] = 8'hc8;
  assign lookUpTable[8'hb2] = 8'h37;
  assign lookUpTable[8'hb3] = 8'h6d;
  assign lookUpTable[8'hb4] = 8'h8d;
  assign lookUpTable[8'hb5] = 8'hd5;
  assign lookUpTable[8'hb6] = 8'h4e;
  assign lookUpTable[8'hb7] = 8'ha9;
  assign lookUpTable[8'hb8] = 8'h6c;
  assign lookUpTable[8'hb9] = 8'h56;
  assign lookUpTable[8'hba] = 8'hf4;
  assign lookUpTable[8'hbb] = 8'hea;
  assign lookUpTable[8'hbc] = 8'h65;
  assign lookUpTable[8'hbd] = 8'h7a;
  assign lookUpTable[8'hbe] = 8'hae;
  assign lookUpTable[8'hbf] = 8'h08;
  assign lookUpTable[8'hc0] = 8'hba;
  assign lookUpTable[8'hc1] = 8'h78;
  assign lookUpTable[8'hc2] = 8'h25;
  assign lookUpTable[8'hc3] = 8'h2e;
  assign lookUpTable[8'hc4] = 8'h1c;
  assign lookUpTable[8'hc5] = 8'ha6;
  assign lookUpTable[8'hc6] = 8'hb4;
  assign lookUpTable[8'hc7] = 8'hc6;
  assign lookUpTable[8'hc8] = 8'he8;
  assign lookUpTable[8'hc9] = 8'hdd;
  assign lookUpTable[8'hca] = 8'h74;
  assign lookUpTable[8'hcb] = 8'h1f;
  assign lookUpTable[8'hcc] = 8'h4b;
  assign lookUpTable[8'hcd] = 8'hbd;
  assign lookUpTable[8'hce] = 8'h8b;
  assign lookUpTable[8'hcf] = 8'h8a;
  assign lookUpTable[8'hd0] = 8'h70;
  assign lookUpTable[8'hd1] = 8'h3e;
  assign lookUpTable[8'hd2] = 8'hb5;
  assign lookUpTable[8'hd3] = 8'h66;
  assign lookUpTable[8'hd4] = 8'h48;
  assign lookUpTable[8'hd5] = 8'h03;
  assign lookUpTable[8'hd6] = 8'hf6;
  assign lookUpTable[8'hd7] = 8'h0e;
  assign lookUpTable[8'hd8] = 8'h61;
  assign lookUpTable[8'hd9] = 8'h35;
  assign lookUpTable[8'hda] = 8'h57;
  assign lookUpTable[8'hdb] = 8'hb9;
  assign lookUpTable[8'hdc] = 8'h86;
  assign lookUpTable[8'hdd] = 8'hc1;
  assign lookUpTable[8'hde] = 8'h1d;
  assign lookUpTable[8'hdf] = 8'h9e;
  assign lookUpTable[8'he0] = 8'he1;
  assign lookUpTable[8'he1] = 8'hf8;
  assign lookUpTable[8'he2] = 8'h98;
  assign lookUpTable[8'he3] = 8'h11;
  assign lookUpTable[8'he4] = 8'h69;
  assign lookUpTable[8'he5] = 8'hd9;
  assign lookUpTable[8'he6] = 8'h8e;
  assign lookUpTable[8'he7] = 8'h94;
  assign lookUpTable[8'he8] = 8'h9b;
  assign lookUpTable[8'he9] = 8'h1e;
  assign lookUpTable[8'hea] = 8'h87;
  assign lookUpTable[8'heb] = 8'he9;
  assign lookUpTable[8'hec] = 8'hce;
  assign lookUpTable[8'hed] = 8'h55;
  assign lookUpTable[8'hee] = 8'h28;
  assign lookUpTable[8'hef] = 8'hdf;
  assign lookUpTable[8'hf0] = 8'h8c;
  assign lookUpTable[8'hf1] = 8'ha1;
  assign lookUpTable[8'hf2] = 8'h89;
  assign lookUpTable[8'hf3] = 8'h0d;
  assign lookUpTable[8'hf4] = 8'hbf;
  assign lookUpTable[8'hf5] = 8'he6;
  assign lookUpTable[8'hf6] = 8'h42;
  assign lookUpTable[8'hf7] = 8'h68;
  assign lookUpTable[8'hf8] = 8'h41;
  assign lookUpTable[8'hf9] = 8'h99;
  assign lookUpTable[8'hfa] = 8'h2d;
  assign lookUpTable[8'hfb] = 8'h0f;
  assign lookUpTable[8'hfc] = 8'hb0;
  assign lookUpTable[8'hfd] = 8'h54;
  assign lookUpTable[8'hfe] = 8'hbb;
  assign lookUpTable[8'hff] = 8'h16;

endmodule 